`default_nettype none


module Control_Unit(
    input logic start,
    input logic reset,
    input logic
);



endmodule